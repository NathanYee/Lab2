// Tests the finite-state machine, the shift register, and maybe some other things

`include "fsm2.v"
`include "shiftregister.v"
`include "datamemory.v"
`include "addresslatch.v"

`define TICK clk = 1; #10; clk = 0; #10; clk = 1; #10; clk = 0; #10; clk = 1; #10; clk = 0; #10;

module testfsm();
	reg clk, sck, cs, mosi, miso;
	wire miso_we, dm_we, sr_we, addr_we;
	wire [7:0] dm_out, sr_contents;
	wire [6:0] dm_addr;

	// finiteStateMachine fsm(sck, cs, mosi, miso_we, dm_we, addr_we, sr_we);
	fsm2 fsm(clk, sck, cs, mosi, miso_we, dm_we, addr_we, sr_we);
	shiftregister sr(clk, sck, sr_we, dm_out, mosi, sr_contents, miso);
	addresslatch al(clk, sr_contents[6:0], addr_we, dm_addr);
	datamemory dm(clk, dm_out, dm_addr, dm_we, sr_contents);

	initial begin
		$dumpfile("fsm.vcd");
		$dumpvars(0, fsm, sr, al, dm);

		clk = 0; sck = 0; cs = 1; mosi = 0; `TICK;

		cs = 0; `TICK;  // Set chip-select low 

		sck = 0; mosi = 0; `TICK; sck = 1; `TICK; // The address
		sck = 0; mosi = 1; `TICK; sck = 1; `TICK;
		sck = 0; mosi = 0; `TICK; sck = 1; `TICK;
		sck = 0; mosi = 1; `TICK; sck = 1; `TICK;
		sck = 0; mosi = 0; `TICK; sck = 1; `TICK;
		sck = 0; mosi = 1; `TICK; sck = 1; `TICK;
		sck = 0; mosi = 0; `TICK; sck = 1; `TICK;

		sck = 0; mosi = 1; `TICK; sck = 1; `TICK; // Write mode

		sck = 0; mosi = 0; `TICK; sck = 1; `TICK; // Data to write
		sck = 0; mosi = 1; `TICK; sck = 1; `TICK;
		sck = 0; mosi = 0; `TICK; sck = 1; `TICK;
		sck = 0; mosi = 1; `TICK; sck = 1; `TICK;
		sck = 0; mosi = 0; `TICK; sck = 1; `TICK;
		sck = 0; mosi = 1; `TICK; sck = 1; `TICK;
		sck = 0; mosi = 0; `TICK; sck = 1; `TICK;
		sck = 0; mosi = 1; `TICK; sck = 1; `TICK;

		cs = 1; `TICK; cs = 0; `TICK;


		sck = 0; mosi = 0; `TICK; sck = 1; `TICK; // The address
		sck = 0; mosi = 1; `TICK; sck = 1; `TICK;
		sck = 0; mosi = 0; `TICK; sck = 1; `TICK;
		sck = 0; mosi = 1; `TICK; sck = 1; `TICK;
		sck = 0; mosi = 0; `TICK; sck = 1; `TICK;
		sck = 0; mosi = 1; `TICK; sck = 1; `TICK;
		sck = 0; mosi = 0; `TICK; sck = 1; `TICK;

		sck = 0; mosi = 0; `TICK; sck = 1; `TICK; // Read mode

		sck = 0; `TICK; sck = 1; `TICK; // Read the data
		sck = 0; `TICK; sck = 1; `TICK;
		sck = 0; `TICK; sck = 1; `TICK;
		sck = 0; `TICK; sck = 1; `TICK;
		sck = 0; `TICK; sck = 1; `TICK;
		sck = 0; `TICK; sck = 1; `TICK;
		sck = 0; `TICK; sck = 1; `TICK;
		sck = 0; `TICK; sck = 1; `TICK;

		$finish;
	end
endmodule
