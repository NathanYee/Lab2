//------------------------------------------------------------------------
// Midpoint Check In
//    1) The parallel data input of the shift register is tied to a constant value
//    2) The load is triggered when button 0 is pressed
//    3) Switches 0 and 1 allow manual control of the serial input
//    4) LEDs show the state of the shift register
//------------------------------------------------------------------------

`include "inputconditioner.v"
`include "shiftregister.v"

module midpoint();

endmodule